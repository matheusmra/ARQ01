module Guia_0204;
    reg [7:0]  b1  = 8'b10110100;
    reg [12:0] b2  = 13'b010111000010; 
    reg [9:0]  b3  = 10'b1110111010;  
    reg [15:0] b4  = 16'b110000010011001;
    reg [15:0] b5  = 16'b1011101001011110; 
    reg [3:0]  b41 = 4'o30;  
    reg [3:0]  b51 = 4'hB;  

    // Actions
    initial
        begin : main
        $display ( "a =  0.%8b (2)            ", b1[7:0]); // a.) 0.10110100(2)
        $display("b = 0.%o%o%o%o%o%o (4)", b2[12:11], b2[10:9], b2[8:7], b2[6:5], b2[4:3], b2[2:1]);
        $display ( "c =  0.%10b (2)           ", b3[9:0]); // c.) 0.1110111010(2)
        $display ( "d =  %o.%o%o%o%o%o (4)        ", b41[3:2], b41[1:0], b4[15:14], b4[13:12], b4[11:10], b4[9:8]); // d.) 30.103211(4)
        $display ( "e =  %o%o.%o%o%o%o%o%o (4)    ", b51[3:2], b51[1:0], b5[15:14], b5[13:12], b5[11:10], b5[9:8], b5[7:6], b5[5:4]); // e.) 23.221132(4)
        
        end // main
endmodule // Guia_0204
